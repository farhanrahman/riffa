LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

PACKAGE project_pak IS

CONSTANT clk_per : time := 8 ns;

END PACKAGE project_pak;