LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY test_core IS

END test_core;

ARCHITECTURE synth OF test_core IS
BEGIN

END ARCHITECTURE synth;
